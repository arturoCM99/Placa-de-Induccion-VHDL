library verilog;
use verilog.vl_types.all;
entity Potencia_vlg_vec_tst is
end Potencia_vlg_vec_tst;
