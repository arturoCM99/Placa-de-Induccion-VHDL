library verilog;
use verilog.vl_types.all;
entity PlacaDeInduccion_vlg_vec_tst is
end PlacaDeInduccion_vlg_vec_tst;
