library verilog;
use verilog.vl_types.all;
entity Tiempo_vlg_sample_tst is
    port(
        K0              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Tiempo_vlg_sample_tst;
