library verilog;
use verilog.vl_types.all;
entity Clasificador_vlg_vec_tst is
end Clasificador_vlg_vec_tst;
