library verilog;
use verilog.vl_types.all;
entity MiniDin_vlg_vec_tst is
end MiniDin_vlg_vec_tst;
