library verilog;
use verilog.vl_types.all;
entity bloquegeneral_vlg_vec_tst is
end bloquegeneral_vlg_vec_tst;
