library verilog;
use verilog.vl_types.all;
entity Tiempo_vlg_vec_tst is
end Tiempo_vlg_vec_tst;
